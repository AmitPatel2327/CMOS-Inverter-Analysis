** sch_path: /home/ap23_27/CMOS_INV/NMOS_inv.sch
**.subckt NMOS_inv
XM2 Vout Vin GND GND sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 nf=1 ad=0.29 as=0.29 pd=2.58 ps=2.58 nrd=0.29 nrs=0.29 sa=0 sb=0 sd=0
+ mult=1 m=1
R1 Vdd Vout 1k m=1
C1 Vout 0 4f m=1
V1 Vin GND Pulse(0 5.0 0 500ps 500ps 4ns 10ns 5)
V2 Vdd GND 5
**** begin user architecture code

.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 100ps 30ns
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
